library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

package pack is
	constant Nbits_dac  : integer := 5;
	constant Nbits_symb : integer :=4;
end pack;
