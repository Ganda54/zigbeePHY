library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

-----------------------------------------------
--zigbee package
--Authors: A & S Ouedraogo
-----------------------------------------------
package pack is
	constant Nbits_dac  : integer := 5;
	constant Nbits_symb : integer :=4;
end pack;
